IceboardTest_SimpleReadWrite2.v