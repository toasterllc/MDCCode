initial begin : test
CLK     <=  1'b0;
CKE     <=  1'b0;
CS_N    <=  1'bz;
RAS_N   <=  1'bz;
CAS_N   <=  1'bz;
WE_N    <=  1'bz;
DM      <=  {DM_BITS{1'bz}};   
ADDR    <=  {ADDR_BITS{1'bz}}; 
BA      <=  2'bzz;			    
Dq      <=  {DQ_BITS  {1'bz}}; 
power_up(200000);
precharge('h00000000, 1);
nop(trp);
refresh;
nop(trfc);
refresh;
nop(trfc);
load_mode('h0, 'h00000033);
nop(tmrd-1);
load_mode('h2, 'h00002000);
nop(tmrd-1);
nop('h000000C8);
activate('h00000000, 'h00000000);
nop(trcd-1);
write(1'b1, 'h00000000, 'h00000004, 1'b1, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0008, 16'h0007, 16'h0006, 16'h0005, 16'h0004, 16'h0003, 16'h0002, 16'h0001});
nop('h00000014);
activate('h00000001, 'h00000000);
nop(trcd-1);
write(1'b1, 'h00000001, 'h00000004, 1'b1, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0018, 16'h0017, 16'h0016, 16'h0015, 16'h0014, 16'h0013, 16'h0012, 16'h0011});
nop('h00000014);
activate('h00000002, 'h00000000);
nop(trcd-1);
write(1'b1, 'h00000002, 'h00000004, 1'b1, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0028, 16'h0027, 16'h0026, 16'h0025, 16'h0024, 16'h0023, 16'h0022, 16'h0021});
nop('h00000014);
activate('h00000003, 'h00000000);
nop(trcd-1);
write(1'b1, 'h00000003, 'h00000004, 1'b1, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0038, 16'h0037, 16'h0036, 16'h0035, 16'h0034, 16'h0033, 16'h0032, 16'h0031});
nop('h00000014);
activate('h00000000, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000000, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0008, 16'h0007, 16'h0006, 16'h0005, 16'h0004, 16'h0003, 16'h0002, 16'h0001});
nop(tras-trcd-1);
precharge('h00000000, 0);
nop('h00000009);
activate('h00000000, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000000, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0008, 16'h0007, 16'h0006, 16'h0005, 16'h0004, 16'h0003, 16'h0002, 16'h0001});
nop(tras-trcd-1);
precharge('h00000000, 0);
nop('h00000009);
activate('h00000000, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000000, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0008, 16'h0007, 16'h0006, 16'h0005, 16'h0004, 16'h0003, 16'h0002, 16'h0001});
nop(tras-trcd-1);
precharge('h00000000, 0);
nop('h00000009);
activate('h00000000, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000000, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0008, 16'h0007, 16'h0006, 16'h0005, 16'h0004, 16'h0003, 16'h0002, 16'h0001});
nop(tras-trcd-1);
precharge('h00000000, 0);
nop('h00000009);
activate('h00000000, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000000, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0008, 16'h0007, 16'h0006, 16'h0005, 16'h0004, 16'h0003, 16'h0002, 16'h0001});
nop(tras-trcd-1);
precharge('h00000000, 0);
nop('h00000009);
activate('h00000000, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000000, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0008, 16'h0007, 16'h0006, 16'h0005, 16'h0004, 16'h0003, 16'h0002, 16'h0001});
nop(tras-trcd-1);
precharge('h00000000, 0);
nop('h00000009);
activate('h00000000, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000000, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0008, 16'h0007, 16'h0006, 16'h0005, 16'h0004, 16'h0003, 16'h0002, 16'h0001});
nop(tras-trcd-1);
precharge('h00000000, 0);
nop('h00000009);
activate('h00000000, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000000, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0008, 16'h0007, 16'h0006, 16'h0005, 16'h0004, 16'h0003, 16'h0002, 16'h0001});
nop(tras-trcd-1);
precharge('h00000000, 0);
nop('h00000009);
activate('h00000000, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000000, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0008, 16'h0007, 16'h0006, 16'h0005, 16'h0004, 16'h0003, 16'h0002, 16'h0001});
nop(tras-trcd-1);
precharge('h00000000, 0);
activate('h00000001, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000001, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0018, 16'h0017, 16'h0016, 16'h0015, 16'h0014, 16'h0013, 16'h0012, 16'h0011});
nop(tras-trcd-1);
precharge('h00000001, 0);
nop('h00000009);
activate('h00000001, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000001, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0018, 16'h0017, 16'h0016, 16'h0015, 16'h0014, 16'h0013, 16'h0012, 16'h0011});
nop(tras-trcd-1);
precharge('h00000001, 0);
nop('h00000009);
activate('h00000001, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000001, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0018, 16'h0017, 16'h0016, 16'h0015, 16'h0014, 16'h0013, 16'h0012, 16'h0011});
nop(tras-trcd-1);
precharge('h00000001, 0);
nop('h00000009);
activate('h00000001, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000001, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0018, 16'h0017, 16'h0016, 16'h0015, 16'h0014, 16'h0013, 16'h0012, 16'h0011});
nop(tras-trcd-1);
precharge('h00000001, 0);
nop('h00000009);
activate('h00000001, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000001, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0018, 16'h0017, 16'h0016, 16'h0015, 16'h0014, 16'h0013, 16'h0012, 16'h0011});
nop(tras-trcd-1);
precharge('h00000001, 0);
nop('h00000009);
activate('h00000001, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000001, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0018, 16'h0017, 16'h0016, 16'h0015, 16'h0014, 16'h0013, 16'h0012, 16'h0011});
nop(tras-trcd-1);
precharge('h00000001, 0);
nop('h00000009);
activate('h00000001, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000001, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0018, 16'h0017, 16'h0016, 16'h0015, 16'h0014, 16'h0013, 16'h0012, 16'h0011});
nop(tras-trcd-1);
precharge('h00000001, 0);
nop('h00000009);
activate('h00000001, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000001, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0018, 16'h0017, 16'h0016, 16'h0015, 16'h0014, 16'h0013, 16'h0012, 16'h0011});
nop(tras-trcd-1);
precharge('h00000001, 0);
nop('h00000009);
activate('h00000001, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000001, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0018, 16'h0017, 16'h0016, 16'h0015, 16'h0014, 16'h0013, 16'h0012, 16'h0011});
nop(tras-trcd-1);
precharge('h00000001, 0);
activate('h00000002, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000002, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0028, 16'h0027, 16'h0026, 16'h0025, 16'h0024, 16'h0023, 16'h0022, 16'h0021});
nop(tras-trcd-1);
precharge('h00000002, 0);
nop('h00000009);
activate('h00000002, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000002, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0028, 16'h0027, 16'h0026, 16'h0025, 16'h0024, 16'h0023, 16'h0022, 16'h0021});
nop(tras-trcd-1);
precharge('h00000002, 0);
nop('h00000009);
activate('h00000002, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000002, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0028, 16'h0027, 16'h0026, 16'h0025, 16'h0024, 16'h0023, 16'h0022, 16'h0021});
nop(tras-trcd-1);
precharge('h00000002, 0);
nop('h00000009);
activate('h00000002, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000002, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0028, 16'h0027, 16'h0026, 16'h0025, 16'h0024, 16'h0023, 16'h0022, 16'h0021});
nop(tras-trcd-1);
precharge('h00000002, 0);
nop('h00000009);
activate('h00000002, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000002, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0028, 16'h0027, 16'h0026, 16'h0025, 16'h0024, 16'h0023, 16'h0022, 16'h0021});
nop(tras-trcd-1);
precharge('h00000002, 0);
nop('h00000009);
activate('h00000002, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000002, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0028, 16'h0027, 16'h0026, 16'h0025, 16'h0024, 16'h0023, 16'h0022, 16'h0021});
nop(tras-trcd-1);
precharge('h00000002, 0);
nop('h00000009);
activate('h00000002, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000002, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0028, 16'h0027, 16'h0026, 16'h0025, 16'h0024, 16'h0023, 16'h0022, 16'h0021});
nop(tras-trcd-1);
precharge('h00000002, 0);
nop('h00000009);
activate('h00000002, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000002, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0028, 16'h0027, 16'h0026, 16'h0025, 16'h0024, 16'h0023, 16'h0022, 16'h0021});
nop(tras-trcd-1);
precharge('h00000002, 0);
nop('h00000009);
activate('h00000002, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000002, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0028, 16'h0027, 16'h0026, 16'h0025, 16'h0024, 16'h0023, 16'h0022, 16'h0021});
nop(tras-trcd-1);
precharge('h00000002, 0);
nop('h00000009);
activate('h00000003, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000003, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0038, 16'h0037, 16'h0036, 16'h0035, 16'h0034, 16'h0033, 16'h0032, 16'h0031});
nop(tras-trcd-1);
precharge('h00000003, 0);
nop('h00000009);
activate('h00000003, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000003, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0038, 16'h0037, 16'h0036, 16'h0035, 16'h0034, 16'h0033, 16'h0032, 16'h0031});
nop(tras-trcd-1);
precharge('h00000003, 0);
nop('h00000009);
activate('h00000003, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000003, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0038, 16'h0037, 16'h0036, 16'h0035, 16'h0034, 16'h0033, 16'h0032, 16'h0031});
nop(tras-trcd-1);
precharge('h00000003, 0);
nop('h00000009);
activate('h00000003, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000003, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0038, 16'h0037, 16'h0036, 16'h0035, 16'h0034, 16'h0033, 16'h0032, 16'h0031});
nop(tras-trcd-1);
precharge('h00000003, 0);
nop('h00000009);
activate('h00000003, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000003, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0038, 16'h0037, 16'h0036, 16'h0035, 16'h0034, 16'h0033, 16'h0032, 16'h0031});
nop(tras-trcd-1);
precharge('h00000003, 0);
nop('h00000009);
activate('h00000003, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000003, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0038, 16'h0037, 16'h0036, 16'h0035, 16'h0034, 16'h0033, 16'h0032, 16'h0031});
nop(tras-trcd-1);
precharge('h00000003, 0);
nop('h00000009);
activate('h00000003, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000003, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0038, 16'h0037, 16'h0036, 16'h0035, 16'h0034, 16'h0033, 16'h0032, 16'h0031});
nop(tras-trcd-1);
precharge('h00000003, 0);
nop('h00000009);
activate('h00000003, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000003, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0038, 16'h0037, 16'h0036, 16'h0035, 16'h0034, 16'h0033, 16'h0032, 16'h0031});
nop(tras-trcd-1);
precharge('h00000003, 0);
nop('h00000009);
activate('h00000003, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000003, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0038, 16'h0037, 16'h0036, 16'h0035, 16'h0034, 16'h0033, 16'h0032, 16'h0031});
nop(tras-trcd-1);
precharge('h00000003, 0);
nop('h00000009);
activate('h00000000, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000000, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0008, 16'h0007, 16'h0006, 16'h0005, 16'h0004, 16'h0003, 16'h0002, 16'h0001});
nop(tras-trcd-1);
precharge('h00000000, 0);
activate('h00000001, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000001, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0018, 16'h0017, 16'h0016, 16'h0015, 16'h0014, 16'h0013, 16'h0012, 16'h0011});
nop(tras-trcd-1);
precharge('h00000001, 0);
activate('h00000002, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000002, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0028, 16'h0027, 16'h0026, 16'h0025, 16'h0024, 16'h0023, 16'h0022, 16'h0021});
nop(tras-trcd-1);
precharge('h00000002, 0);
activate('h00000003, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000003, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0038, 16'h0037, 16'h0036, 16'h0035, 16'h0034, 16'h0033, 16'h0032, 16'h0031});
nop(tras-trcd-1);
precharge('h00000003, 0);
activate('h00000000, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000000, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0008, 16'h0007, 16'h0006, 16'h0005, 16'h0004, 16'h0003, 16'h0002, 16'h0001});
nop(tras-trcd-1);
precharge('h00000000, 0);
activate('h00000001, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000001, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0018, 16'h0017, 16'h0016, 16'h0015, 16'h0014, 16'h0013, 16'h0012, 16'h0011});
nop(tras-trcd-1);
precharge('h00000001, 0);
activate('h00000002, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000002, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0028, 16'h0027, 16'h0026, 16'h0025, 16'h0024, 16'h0023, 16'h0022, 16'h0021});
nop(tras-trcd-1);
precharge('h00000002, 0);
activate('h00000003, 'h00000000);
nop(trcd-1);
read_verify(1'b1, 'h00000003, 'h00000004, 1'b0, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0}, {16'h0038, 16'h0037, 16'h0036, 16'h0035, 16'h0034, 16'h0033, 16'h0032, 16'h0031});
nop(tras-trcd-1);
precharge('h00000003, 0);
nop('h0000000A);
test_done;
end


