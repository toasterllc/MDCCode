IcestickSDRAMTest.v