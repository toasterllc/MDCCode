Top.v