IcestickTest_SDRAMReadWriteRandomly.v