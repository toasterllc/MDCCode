IceboardTest_SDRAMReadWriteRandomly.v