`define SYNTH
`include "SDRAMController.v"

module Top();
endmodule
