`timescale 1ns/1ps
`include "../ClockGen.v"
`include "../SDRAMController.v"
`include "../uart.v"

`ifdef SIM
`include "../mt48h32m16lf/mobile_sdr.v"
`endif

module Top(
    input wire          clk12mhz,
    
    output wire[7:0]    led,
    
    output wire         ram_clk,
    output wire         ram_cke,
    output wire[1:0]    ram_ba,
    output wire[12:0]   ram_a,
    output wire         ram_cs_,
    output wire         ram_ras_,
    output wire         ram_cas_,
    output wire         ram_we_,
    output wire[1:0]    ram_dqm,
    inout wire[15:0]    ram_dq,
    
    input wire          uart_rx,
    output wire         uart_tx
);
    function [15:0] DataFromAddr;
        input [24:0] addr;
        // DataFromAddr = {7'h55, addr[24:16]} ^ ~(addr[15:0]);
        DataFromAddr = addr[15:0];
        // DataFromAddr = 16'hFFFF;
        // DataFromAddr = 16'h0000;
        // DataFromAddr = 16'h7832;
    endfunction
    
    // 24 MHz clock
    localparam ClockFrequency = 24000000;
    wire clk;
    wire rst;
    ClockGen #(
        .FREQ(ClockFrequency),
		.DIVR(0),
		.DIVF(63),
		.DIVQ(5),
		.FILTER_RANGE(1)
    ) cg(.clk12mhz(clk12mhz), .clk(clk), .rst(rst));
    
    localparam AddrWidth = 25;
    localparam AddrCount = 'h2000000;
    localparam AddrCountLimit = AddrCount;
    // localparam AddrCountLimit = 'h10000;
    // localparam AddrCountLimit = AddrCount/8192;
    
    
    // localparam AddrCountLimit = AddrCount/512;
    // localparam AddrCountLimit = AddrCount/1024; // 32k words
    // localparam AddrCountLimit = AddrCount/8192;
    localparam DataWidth = 16;
    
    localparam StatusStart          = 0;
    localparam StatusInit           = 1;
    localparam StatusUnderway       = 2;
    localparam StatusTooManyReads   = 3;
    localparam StatusInvalidData    = 4;
    localparam StatusUnexpectedData = 5;
    
    wire                  cmdReady;
    reg                   cmdTrigger = 0;
    reg[AddrWidth-1:0]    cmdAddr = 0;
    reg                   cmdWrite = 0;
    reg[DataWidth-1:0]    cmdWriteData = 0;
    wire[DataWidth-1:0]   cmdReadData;
    wire                  cmdReadDataValid;
    
    localparam MaxEnqueuedReads = 10;
    reg[(AddrWidth*MaxEnqueuedReads)-1:0] readAddr = 0;
    reg[$clog2(MaxEnqueuedReads)-1:0] enqueuedReadCount = 0;
    
    wire[AddrWidth-1:0] currentReadAddr = readAddr[AddrWidth-1:0];
    wire[DataWidth-1:0] expectedReadData = DataFromAddr(currentReadAddr);
    
    reg[6:0] status = StatusStart /* synthesis syn_keep=1 */; // syn_keep is necessary to prevent Synplify optimization from removing -- "removing sequential instance ..."
    assign led[6:0] = status;
    
    reg wrapped = 0;
    assign led[7] = wrapped;
    
    SDRAMController #(
        .ClockFrequency(ClockFrequency)
    ) sdramController(
        .clk(clk),
        
        .cmdReady(cmdReady),
        .cmdTrigger(cmdTrigger),
        .cmdAddr(cmdAddr),
        .cmdWrite(cmdWrite),
        .cmdWriteData(cmdWriteData),
        .cmdReadData(cmdReadData),
        .cmdReadDataValid(cmdReadDataValid),
        
        .ram_clk(ram_clk),
        .ram_cke(ram_cke),
        .ram_ba(ram_ba),
        .ram_a(ram_a),
        .ram_cs_(ram_cs_),
        .ram_ras_(ram_ras_),
        .ram_cas_(ram_cas_),
        .ram_we_(ram_we_),
        .ram_dqm(ram_dqm),
        .ram_dq(ram_dq)
    );
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    // UART stuff
    reg uartTransmit = 0;
    reg [7:0] uartTxByte = 0;
    wire uartReceived;
    wire [7:0] uartRxByte;
    wire uartReceiving;
    wire uartTransmitting;
    
    uart #(
        .baud_rate(9600),                   // The baud rate in kilobits/s
        .sys_clk_freq(ClockFrequency)       // The master clock frequency
    )
    uart0(
        .clk(clk),                          // The master clock for this module
        .rst(rst),                          // Synchronous reset
        .rx(uart_rx),                       // Incoming serial line
        .tx(uart_tx),                       // Outgoing serial line
        .transmit(uartTransmit),            // Signal to transmit
        .tx_byte(uartTxByte),               // Byte to transmit
        .received(uartReceived),            // Indicated that a byte has been received
        .rx_byte(uartRxByte),               // Byte received
        .is_receiving(uartReceiving),       // Low when receive line is idle
        .is_transmitting(uartTransmitting), // Low when transmit line is idle
        .recv_error()                       // Indicates error in receiving packet.
    );
    
    reg[2:0]      uartStage = 0;
    
    reg[63:0]     uartDataIn = 0;
    reg[15:0]     uartDataInCount = 0;
    reg           uartDataInSuppress = 0;
    
    reg[32*8-1:0] uartDataOut = 0;
    reg[15:0]     uartDataOutCount = 0;
    
    function [7:0] HexASCIIFromNibble;
        input [3:0] n;
        HexASCIIFromNibble = (n<10 ? 8'd48+n : 8'd97-8'd10+n);
    endfunction
    
    function [3:0] NibbleFromHexASCII;
        input [7:0] n;
        NibbleFromHexASCII = (n>=97 ? n-97+10 : n-48);
    endfunction
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    task Read(input [AddrWidth-1:0] addr); begin
        cmdTrigger <= 1;
        cmdAddr <= addr;
        cmdWrite <= 0;
        
        if (enqueuedReadCount >= MaxEnqueuedReads) begin
            `ifdef SIM
                $error("Too many enqueued reads");
            `endif
            
            status <= StatusTooManyReads;
        end
        
        readAddr <= (addr<<(AddrWidth*enqueuedReadCount))|readAddr;
        enqueuedReadCount <= enqueuedReadCount+1;
    end endtask
    
    always @(posedge clk) begin
        // Set our default state if the current command was accepted
        if (cmdReady) cmdTrigger <= 0;
        
        // By default we're not transmitting
        uartTransmit <= 0;
        
        // Transmit another UART byte if data is available, and we're not currently transmitting
        if (!uartTransmit && !uartTransmitting && uartDataOutCount>0) begin
			uartTxByte <= uartDataOut[(8*uartDataOutCount)-1 -: 8];
            uartTransmit <= 1;
			uartDataOutCount <= uartDataOutCount-1;
        end
        
        // Initialize memory to known values
        if (status == StatusStart) begin
            cmdTrigger <= 1;
            cmdAddr <= 0;
            cmdWrite <= 1;
            cmdWriteData <= DataFromAddr(0);
            
            status <= StatusInit;
        
        end else if (status == StatusInit) begin
            // The SDRAM controller accepted the command, so transition to the next state
            if (cmdReady) begin
                if (cmdAddr < AddrCountLimit-1) begin
                    cmdTrigger <= 1;
                    cmdAddr <= cmdAddr+1;
                    cmdWrite <= 1;
                    cmdWriteData <= DataFromAddr(cmdAddr+1);
                    
                    `ifdef SIM
                        if (!(cmdAddr % 'h1000)) begin
                            $display("Initializing memory: %h", cmdAddr);
                        end
                    `endif
                
                end else begin
                    // Kick off reading
                    Read(0);
                    
                    // Next stage
                    status <= StatusUnderway;
                end
                
                // $display("Write: %h", cmdAddr);
            end
        
        end else begin
            // Handle read data if available
            if (cmdReadDataValid) begin
                if (enqueuedReadCount > 0) begin
                    // $display("Read data: 0x%h", cmdReadData);
                    
                    // Verify that the data read out is what we expect
                    if (cmdReadData != expectedReadData) begin
                        `ifdef SIM
                            $error("Read invalid data (expected: 0x%h, got: 0x%h)", expectedReadData, cmdReadData);
                        `endif
                        
                        status <= StatusInvalidData;
                        
                        if (uartDataOutCount == 0) begin
                            uartDataOut <= {
                                HexASCIIFromNibble({3'b0, currentReadAddr[24:24]}),
                                HexASCIIFromNibble(currentReadAddr[23:20]),
                                HexASCIIFromNibble(currentReadAddr[19:16]),
                                HexASCIIFromNibble(currentReadAddr[15:12]),
                                HexASCIIFromNibble(currentReadAddr[11:8]),
                                HexASCIIFromNibble(currentReadAddr[7:4]),
                                HexASCIIFromNibble(currentReadAddr[3:0]),
                            
                                "E",
                                HexASCIIFromNibble(expectedReadData[15:12]),
                                HexASCIIFromNibble(expectedReadData[11:8]),
                                HexASCIIFromNibble(expectedReadData[7:4]),
                                HexASCIIFromNibble(expectedReadData[3:0]),
                            
                                "G",
                                HexASCIIFromNibble(cmdReadData[15:12]),
                                HexASCIIFromNibble(cmdReadData[11:8]),
                                HexASCIIFromNibble(cmdReadData[7:4]),
                                HexASCIIFromNibble(cmdReadData[3:0]),
                            
                                "\r\n"
                            };
                            
                            uartDataOutCount <= 19;
                        end
                        
                    end else begin
                        $display("Read expected data from addr 0x%x: 0x%x", currentReadAddr, DataFromAddr(currentReadAddr));
                    end
                    
                    readAddr <= readAddr >> AddrWidth;
                    enqueuedReadCount <= enqueuedReadCount-1;
                
                // Something's wrong if we weren't expecting data and we got some
                end else begin
                    `ifdef SIM
                        $error("Received data when we didn't expect any");
                    `endif
                    
                    status <= StatusUnexpectedData;
                end
            end
            
            // Current command was accepted: prepare a new command
            else if (cmdReady) begin
                // A command was accepted, issue a new one
                // `ifdef SIM
                //     $display("Enqueue read @ 0x%h", cmdAddr);
                // `endif
                
                Read((cmdAddr+1)&(AddrCountLimit-1));
                
                if (cmdAddr == 0) begin
                    wrapped <= !wrapped;
                end
            end
        end
    end
    
`ifdef SIM
    mobile_sdr sdram(
        .clk(ram_clk),
        .cke(ram_cke),
        .addr(ram_a),
        .ba(ram_ba),
        .cs_n(ram_cs_),
        .ras_n(ram_ras_),
        .cas_n(ram_cas_),
        .we_n(ram_we_),
        .dq(ram_dq),
        .dqm(ram_dqm)
    );
    
    // initial begin
    //     $dumpfile("top.vcd");
    //     $dumpvars(0, Top);
    //     // #1000000000;
    //     // $finish;
    // end
`endif
endmodule
