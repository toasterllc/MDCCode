blink.v