`include "Util.v"
`include "ClockGen.v"
`include "AFIFO.v"
`include "ToggleAck.v"
`include "TogglePulse.v"

`timescale 1ps/1ps

`ifdef SIM
localparam ImageWidth = 2304;
// localparam ImageHeight = 1296;
localparam ImageHeight = 16;
`else
localparam ImageWidth = 6000;
localparam ImageHeight = 6000;
`endif

localparam ImageSize = ImageWidth*ImageHeight;

module Top(
    input wire          clk24mhz,
    output reg[3:0]     led = 0
);
    // ====================
    // Clock (97.5 MHz)
    // ====================
    localparam PixDClkFreq = 97_500_000;
    wire pix_dclk;
    ClockGen #(
        .FREQ(PixDClkFreq),
        .DIVR(1),
        .DIVF(64),
        .DIVQ(3),
        .FILTER_RANGE(1)
    ) ClockGen_pix_dclk(.clkRef(clk24mhz), .clk(pix_dclk));
    
    // ====================
    // Clock (120 MHz)
    // ====================
    localparam ClkFreq = 120_000_000;
    wire clk;
    ClockGen #(
        .FREQ(ClkFreq),
        .DIVR(0),
        .DIVF(39),
        .DIVQ(3),
        .FILTER_RANGE(2)
    ) ClockGen_clk(.clkRef(clk24mhz), .clk(clk));
    
    // ====================
    // FIFO
    // ====================
    reg fifo_writeEn = 0;
    wire fifo_writeReady;
    reg fifo_readTrigger = 0;
    wire[15:0] fifo_readData;
    wire fifo_readReady;
    reg[`RegWidth(ImageSize-1)-1:0] fifo_counter = 0;
        
    AFIFO #(
        .Width(16),
        .Size(256)
    ) AFIFO (
        .wclk(pix_dclk),
        .wok(fifo_writeReady),
        .wtrigger(fifo_writeEn),
        .wdata({3'b0, fifo_counter}),
        
        .rclk(clk),
        .rok(fifo_readReady),
        .rtrigger(fifo_readTrigger),
        .rdata(fifo_readData)
    );
    
    reg ctrl_fifoCaptureTrigger = 0;
    `TogglePulse(fifo_captureTrigger, ctrl_fifoCaptureTrigger, posedge, pix_dclk);
    
    reg[2:0] fifo_state = 0;
    always @(posedge pix_dclk) begin
        fifo_writeEn <= 0; // Reset by default
        
        case (fifo_state)
        // Idle: wait to be triggered
        0: begin
        end
        
        // Wait for FIFO to be done resetting
        1: begin
            $display("[FIFO] Frame start");
            fifo_counter <= ImageSize-1;
            fifo_state <= 2;
        end
        
        // Wait until the end of the frame
        2: begin
            fifo_writeEn <= 1;
            if (fifo_writeEn) begin
                if (fifo_writeReady) begin
                    fifo_counter <= fifo_counter-1;
                    if (!fifo_counter) begin
                        $display("[FIFO] Frame end");
                        fifo_writeEn <= 0;
                        fifo_state <= 0;
                    end
                
                end else begin
                    $display("[FIFO] Pixel dropped ❌");
                    led[2] <= 1;
                    `Finish;
                end
            end
        end
        endcase
        
        if (fifo_captureTrigger) begin
            fifo_state <= 1;
        end
    end
    
    
    
    reg[2:0] ctrl_state = 0;
    reg[`RegWidth(ImageSize-1)-1:0] ctrl_pixelCounter = 0;
    reg[9:0] ctrl_counter = 0;
    always @(posedge clk) begin
        ctrl_counter <= ctrl_counter+1;
        fifo_readTrigger <= 0;
        
        case (ctrl_state)
        0: begin
            if (&ctrl_counter) begin
                ctrl_state <= 1;
            end
        end
        
        1: begin
            $display("[CTRL] Triggered");
            led[0] <= !led[0];
            ctrl_state <= 2;
        end
        
        2: begin
            // Start the FIFO data flow
            ctrl_fifoCaptureTrigger <= !ctrl_fifoCaptureTrigger;
            ctrl_pixelCounter <= ImageSize-1;
            ctrl_state <= 3;
        end
        
        // Receive data out of FIFO
        3: begin
            fifo_readTrigger <= 1;
            
            if (fifo_readTrigger && fifo_readReady) begin
                $display("[CTRL] Got pixel: %0d (%0d)", fifo_readData, ctrl_pixelCounter);
                ctrl_pixelCounter <= ctrl_pixelCounter-1;
                if (!ctrl_pixelCounter) begin
                    $display("[CTRL] Received full image");
                    fifo_readTrigger <= 0;
                    ctrl_state <= 4;
                end
            end
        end
        
        // Wait for extra pixels that we don't expect
        4: begin
            if (fifo_readReady) begin
                // We got a pixel we didn't expect
                $display("[CTRL] Got extra pixel ❌");
                led[3] <= !led[3];
                `Finish;
            end
        end
        endcase
    end
endmodule








`ifdef SIM
module Testbench();
    reg clk24mhz = 0;
    wire[3:0] led;
    
    Top Top(.*);
    
    // initial begin
    //     $dumpfile("Top.vcd");
    //     $dumpvars(0, Testbench);
    // end
endmodule
`endif
