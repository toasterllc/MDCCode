test.v