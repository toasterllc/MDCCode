IceboardTest_Blinky.v