IceboardTest_SDRAMReadWriteViaUART.v