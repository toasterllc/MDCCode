IcestickTest_SDRAMReadWriteViaUART.v