top.v